
module AvalonMM_hyperRamS27KL0641_interface (
	clk_clk,
	reset_reset_n);	

	input		clk_clk;
	input		reset_reset_n;
endmodule
