-- AvalonMM_hyperRamS27KL0641_interface.vhd

-- Generated using ACDS version 22.1 917

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity AvalonMM_hyperRamS27KL0641_interface is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity AvalonMM_hyperRamS27KL0641_interface;

architecture rtl of AvalonMM_hyperRamS27KL0641_interface is
begin

end architecture rtl; -- of AvalonMM_hyperRamS27KL0641_interface
