-- unsaved.vhd

-- Generated using ACDS version 22.1 917

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unsaved is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity unsaved;

architecture rtl of unsaved is
begin

end architecture rtl; -- of unsaved
